LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.numeric_std.ALL;

ENTITY Control_Unit IS
	PORT (
		rst : IN STD_LOGIC;
		opcode : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
		Flag_Enable : OUT STD_LOGIC;
		OutPort_Enable : OUT STD_LOGIC;
		RegWrite : OUT STD_LOGIC;
		Address: OUT STD_LOGIC;
		INT_sig: OUT STD_LOGIC;
		MemRead : OUT STD_LOGIC;
		MemWrite : OUT STD_LOGIC;
		MTR : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
		SP_sig : OUT STD_LOGIC_VECTOR (1 DOWNTO 0); -- SP[1] = PLUS; SP[0] = MINUS
		FR: OUT STD_LOGIC;
		Write_Data_sel : OUT STD_LOGIC;
		RET_sig: OUT STD_LOGIC;
		JZ: OUT STD_LOGIC;
		JN: OUT STD_LOGIC;
		JC: OUT STD_LOGIC;
		ALU_sel : OUT STD_LOGIC_VECTOR (2 DOWNTO 0);
		JMP_branch : OUT STD_LOGIC;
		UC: OUT STD_LOGIC;
		RdRs_sel: OUT STD_LOGIC;
		Rsrc1_Rscr2_sel : OUT STD_LOGIC;
		PC_disable: OUT STD_LOGIC
	);
END ENTITY Control_Unit;

ARCHITECTURE Control_Unit_arch OF Control_Unit IS
BEGIN
	PROCESS (opcode, rst) IS
	BEGIN
		IF(rst = '1') THEN
			-- Reset all outputs to their default state
			Flag_Enable       <= '0';
			OutPort_Enable    <= '0';
			RegWrite          <= '0';
			Address           <= '0';
			INT_sig           <= '0';
			MemRead           <= '0';
			MemWrite          <= '0';
			MTR               <= (others => '0');
			SP_sig            <= (others => '0');
			FR                <= '0';
			Write_Data_sel    <= '0';
			RET_sig           <= '0';
			JZ                <= '0';
			JN                <= '0';
			JC                <= '0';
			ALU_sel           <= (others => '0');    
			JMP_branch        <= '0';
			UC                <= '0';
			RdRs_sel          <= '0';
			Rsrc1_Rscr2_sel   <= '0';
			PC_disable        <= '0';
      ELSE
			IF (opcode = "00000") THEN --NOP
				Flag_Enable       <= '0';
				OutPort_Enable    <= '0';
				RegWrite          <= '0';
				Address           <= '0';
				INT_sig           <= '0';
				MemRead           <= '0';
				MemWrite          <= '0';
				MTR               <= (others => '0');
				SP_sig            <= (others => '0');
				FR                <= '0';
				Write_Data_sel    <= '0';
				RET_sig           <= '0';
				JZ                <= '0';
				JN                <= '0';
				JC                <= '0';
				ALU_sel           <= "000";
				JMP_branch        <= '0';
				UC                <= '0';
				RdRs_sel          <= '0';
				Rsrc1_Rscr2_sel   <= '0';
				PC_disable        <= '0';
			END IF;
			IF (opcode = "00001") THEN --HLT
				Flag_Enable       <= '0';
				OutPort_Enable    <= '0';
				RegWrite          <= '0';
				Address           <= '0';
				INT_sig           <= '0';
				MemRead           <= '0';
				MemWrite          <= '0';
				MTR               <= (others => '0');
				SP_sig            <= (others => '0');
				FR                <= '0';
				Write_Data_sel    <= '0';
				RET_sig           <= '0';
				JZ                <= '0';
				JN                <= '0';
				JC                <= '0';
				ALU_sel           <= "000";
				JMP_branch        <= '0';
				UC                <= '0';
				RdRs_sel          <= '0';
				Rsrc1_Rscr2_sel   <= '0';
				PC_disable        <= '1';
			END IF;
			IF (opcode = "00010") THEN --SETC
				Flag_Enable       <= '1';
				OutPort_Enable    <= '0';
				RegWrite          <= '0';
				Address           <= '0';
				INT_sig           <= '0';
				MemRead           <= '0';
				MemWrite          <= '0';
				MTR               <= (others => '0');
				SP_sig            <= (others => '0');
				FR                <= '0';
				Write_Data_sel    <= '0';
				RET_sig           <= '0';
				JZ                <= '0';
				JN                <= '0';
				JC                <= '0';
				ALU_sel           <= "011";
				JMP_branch        <= '0';
				UC                <= '0';
				RdRs_sel          <= '0';
				Rsrc1_Rscr2_sel   <= '0';
				PC_disable        <= '0';
			END IF;
			IF (opcode = "00011") THEN --NOT
				Flag_Enable       <= '1';
				OutPort_Enable    <= '0';
				RegWrite          <= '1';
				Address           <= '0';
				INT_sig           <= '0';
				MemRead           <= '0';
				MemWrite          <= '0';
				MTR               <= (others => '0');
				SP_sig            <= (others => '0');
				FR                <= '0';
				Write_Data_sel    <= '0';
				RET_sig           <= '0';
				JZ                <= '0';
				JN                <= '0';
				JC                <= '0';
				ALU_sel           <= "000";
				JMP_branch        <= '0';
				UC                <= '0';
				RdRs_sel          <= '1';
				Rsrc1_Rscr2_sel   <= '0';
				PC_disable        <= '0';
			END IF;
			IF (opcode = "00100") THEN --INC
				Flag_Enable       <= '1';
				OutPort_Enable    <= '0';
				RegWrite          <= '1';
				Address           <= '0';
				INT_sig           <= '0';
				MemRead           <= '0';
				MemWrite          <= '0';
				MTR               <= (others => '0');
				SP_sig            <= (others => '0');
				FR                <= '0';
				Write_Data_sel    <= '0';
				RET_sig           <= '0';
				JZ                <= '0';
				JN                <= '0';
				JC                <= '0';
				ALU_sel           <= "111";
				JMP_branch        <= '0';
				UC                <= '0';
				RdRs_sel          <= '1';
				Rsrc1_Rscr2_sel   <= '0';
				PC_disable        <= '0';
			END IF;
			IF (opcode = "00101") THEN --OUT
				Flag_Enable       <= '0';
				OutPort_Enable    <= '1';
				RegWrite          <= '0';
				Address           <= '0';
				INT_sig           <= '0';
				MemRead           <= '0';
				MemWrite          <= '0';
				MTR               <= (others => '0');
				SP_sig            <= (others => '0');
				FR                <= '0';
				Write_Data_sel    <= '0';
				RET_sig           <= '0';
				JZ                <= '0';
				JN                <= '0';
				JC                <= '0';
				ALU_sel           <= "100";
				JMP_branch        <= '0';
				UC                <= '0';
				RdRs_sel          <= '0';
				Rsrc1_Rscr2_sel   <= '0';
				PC_disable        <= '0';
			END IF;
			IF (opcode = "00110") THEN --IN
				Flag_Enable       <= '0';
				OutPort_Enable    <= '0';
				RegWrite          <= '1';
				Address           <= '0';
				INT_sig           <= '0';
				MemRead           <= '0';
				MemWrite          <= '0';
				MTR               <= "10";
				SP_sig            <= (others => '0');
				FR                <= '0';
				Write_Data_sel    <= '0';
				RET_sig           <= '0';
				JZ                <= '0';
				JN                <= '0';
				JC                <= '0';
				ALU_sel           <= "000";
				JMP_branch        <= '0';
				UC                <= '0';
				RdRs_sel          <= '1';
				Rsrc1_Rscr2_sel   <= '0';
				PC_disable        <= '0';
			END IF;
			IF (opcode = "00111") THEN --MOV
				Flag_Enable       <= '0';
				OutPort_Enable    <= '0';
				RegWrite          <= '1';
				Address           <= '0';
				INT_sig           <= '0';
				MemRead           <= '0';
				MemWrite          <= '0';
				MTR               <= (others => '0');
				SP_sig            <= (others => '0');
				FR                <= '0';
				Write_Data_sel    <= '0';
				RET_sig           <= '0';
				JZ                <= '0';
				JN                <= '0';
				JC                <= '0';
				ALU_sel           <= "100";
				JMP_branch        <= '0';
				UC                <= '0';
				RdRs_sel          <= '1';
				Rsrc1_Rscr2_sel   <= '0';
				PC_disable        <= '0';
			END IF;
			IF (opcode = "01000") THEN --ADD
				Flag_Enable       <= '1';
				OutPort_Enable    <= '0';
				RegWrite          <= '1';
				Address           <= '0';
				INT_sig           <= '0';
				MemRead           <= '0';
				MemWrite          <= '0';
				MTR               <= (others => '0');
				SP_sig            <= (others => '0');
				FR                <= '0';
				Write_Data_sel    <= '0';
				RET_sig           <= '0';
				JZ                <= '0';
				JN                <= '0';
				JC                <= '0';
				ALU_sel           <= "110";
				JMP_branch        <= '0';
				UC                <= '0';
				RdRs_sel          <= '1';
				Rsrc1_Rscr2_sel   <= '0';
				PC_disable        <= '0';
			END IF;
			IF (opcode = "01001") THEN --SUB
				Flag_Enable       <= '1';
				OutPort_Enable    <= '0';
				RegWrite          <= '1';
				Address           <= '0';
				INT_sig           <= '0';
				MemRead           <= '0';
				MemWrite          <= '0';
				MTR               <= (others => '0');
				SP_sig            <= (others => '0');
				FR                <= '0';
				Write_Data_sel    <= '0';
				RET_sig           <= '0';
				JZ                <= '0';
				JN                <= '0';
				JC                <= '0';
				ALU_sel           <= "010";
				JMP_branch        <= '0';
				UC                <= '0';
				RdRs_sel          <= '1';
				Rsrc1_Rscr2_sel   <= '0';
				PC_disable        <= '0';
			END IF;
			IF (opcode = "01010") THEN --AND
				Flag_Enable       <= '1';
				OutPort_Enable    <= '0';
				RegWrite          <= '1';
				Address           <= '0';
				INT_sig           <= '0';
				MemRead           <= '0';
				MemWrite          <= '0';
				MTR               <= (others => '0');
				SP_sig            <= (others => '0');
				FR                <= '0';
				Write_Data_sel    <= '0';
				RET_sig           <= '0';
				JZ                <= '0';
				JN                <= '0';
				JC                <= '0';
				ALU_sel           <= "001";
				JMP_branch        <= '0';
				UC                <= '0';
				RdRs_sel          <= '1';
				Rsrc1_Rscr2_sel   <= '0';
				PC_disable        <= '0';
			END IF;
			IF (opcode = "01011") THEN --IADD
				Flag_Enable       <= '1';
				OutPort_Enable    <= '0';
				RegWrite          <= '1';
				Address           <= '0';
				INT_sig           <= '0';
				MemRead           <= '0';
				MemWrite          <= '0';
				MTR               <= (others => '0');
				SP_sig            <= (others => '0');
				FR                <= '0';
				Write_Data_sel    <= '0';
				RET_sig           <= '0';
				JZ                <= '0';
				JN                <= '0';
				JC                <= '0';
				ALU_sel           <= "110";
				JMP_branch        <= '0';
				UC                <= '0';
				RdRs_sel          <= '1';
				Rsrc1_Rscr2_sel   <= '0';
				PC_disable        <= '0';
			END IF;
			IF (opcode = "01100") THEN --PUSH
				Flag_Enable       <= '0';
				OutPort_Enable    <= '0';
				RegWrite          <= '0';
				Address           <= '1';
				INT_sig           <= '0';
				MemRead           <= '0';
				MemWrite          <= '1';
				MTR               <= "00";
				SP_sig            <= "01";
				FR                <= '0';
				Write_Data_sel    <= '0';
				RET_sig           <= '0';
				JZ                <= '0';
				JN                <= '0';
				JC                <= '0';
				ALU_sel           <= "000";
				JMP_branch        <= '0';
				UC                <= '0';
				RdRs_sel          <= '0';
				Rsrc1_Rscr2_sel   <= '0';
				PC_disable        <= '0';
			END IF;
			IF (opcode = "01101") THEN --POP
				Flag_Enable       <= '0';
				OutPort_Enable    <= '0';
				RegWrite          <= '1';
				Address           <= '1';
				INT_sig           <= '0';
				MemRead           <= '1';
				MemWrite          <= '0';
				MTR               <= "01";
				SP_sig            <= "10";
				FR                <= '0';
				Write_Data_sel    <= '0';
				RET_sig           <= '0';
				JZ                <= '0';
				JN                <= '0';
				JC                <= '0';
				ALU_sel           <= "000";
				JMP_branch        <= '0';
				UC                <= '0';
				RdRs_sel          <= '1';
				Rsrc1_Rscr2_sel   <= '0';
				PC_disable        <= '0';
			END IF;
			IF (opcode = "01110") THEN --LDM
				Flag_Enable       <= '0';
				OutPort_Enable    <= '0';
				RegWrite          <= '1';
				Address           <= '0';
				INT_sig           <= '0';
				MemRead           <= '0';
				MemWrite          <= '0';
				MTR               <= (others => '0');
				SP_sig            <= (others => '0');
				FR                <= '0';
				Write_Data_sel    <= '0';
				RET_sig           <= '0';
				JZ                <= '0';
				JN                <= '0';
				JC                <= '0';
				ALU_sel           <= "101";
				JMP_branch        <= '0';
				UC                <= '0';
				RdRs_sel          <= '1';
				Rsrc1_Rscr2_sel   <= '0';
				PC_disable        <= '0';
			END IF;
			IF (opcode = "01111") THEN --LDD
				Flag_Enable       <= '0';
				OutPort_Enable    <= '0';
				RegWrite          <= '1';
				Address           <= '1';
				INT_sig           <= '0';
				MemRead           <= '1';
				MemWrite          <= '0';
				MTR               <= "01";
				SP_sig            <= (others => '0');
				FR                <= '0';
				Write_Data_sel    <= '0';
				RET_sig           <= '0';
				JZ                <= '0';
				JN                <= '0';
				JC                <= '0';
				ALU_sel           <= "110";
				JMP_branch        <= '0';
				UC                <= '0';
				RdRs_sel          <= '1';
				Rsrc1_Rscr2_sel   <= '0';
				PC_disable        <= '0';
			END IF;
			IF (opcode = "10000") THEN --STD
				Flag_Enable       <= '0';
				OutPort_Enable    <= '0';
				RegWrite          <= '0';
				Address           <= '1';
				INT_sig           <= '0';
				MemRead           <= '0';
				MemWrite          <= '1';
				MTR               <= "00";
				SP_sig            <= (others => '0');
				FR                <= '0';
				Write_Data_sel    <= '0';
				RET_sig           <= '0';
				JZ                <= '0';
				JN                <= '0';
				JC                <= '0';
				ALU_sel           <= "110";
				JMP_branch        <= '0';
				UC                <= '0';
				RdRs_sel          <= '0';
				Rsrc1_Rscr2_sel   <= '1';
				PC_disable        <= '0';
			END IF;
			IF (opcode = "10001") THEN --JZ
				Flag_Enable       <= '0';
				OutPort_Enable    <= '0';
				RegWrite          <= '0';
				Address           <= '0';
				INT_sig           <= '0';
				MemRead           <= '0';
				MemWrite          <= '0';
				MTR               <= "00";
				SP_sig            <= (others => '0');
				FR                <= '0';
				Write_Data_sel    <= '0';
				RET_sig           <= '0';
				JZ                <= '1';
				JN                <= '0';
				JC                <= '0';
				ALU_sel           <= "000";
				JMP_branch        <= '1';
				UC                <= '0';
				RdRs_sel          <= '0';
				Rsrc1_Rscr2_sel   <= '0';
				PC_disable        <= '0';
			END IF;
			IF (opcode = "10010") THEN --JN
				Flag_Enable       <= '0';
				OutPort_Enable    <= '0';
				RegWrite          <= '0';
				Address           <= '0';
				INT_sig           <= '0';
				MemRead           <= '0';
				MemWrite          <= '0';
				MTR               <= "00";
				SP_sig            <= (others => '0');
				FR                <= '0';
				Write_Data_sel    <= '0';
				RET_sig           <= '0';
				JZ                <= '0';
				JN                <= '1';
				JC                <= '0';
				ALU_sel           <= "000";
				JMP_branch        <= '1';
				UC                <= '0';
				RdRs_sel          <= '0';
				Rsrc1_Rscr2_sel   <= '0';
				PC_disable        <= '0';
			END IF;
			IF (opcode = "10011") THEN --JC
				Flag_Enable       <= '0';
				OutPort_Enable    <= '0';
				RegWrite          <= '0';
				Address           <= '0';
				INT_sig           <= '0';
				MemRead           <= '0';
				MemWrite          <= '0';
				MTR               <= "00";
				SP_sig            <= (others => '0');
				FR                <= '0';
				Write_Data_sel    <= '0';
				RET_sig           <= '0';
				JZ                <= '0';
				JN                <= '0';
				JC                <= '1';
				ALU_sel           <= "000";
				JMP_branch        <= '1';
				UC                <= '0';
				RdRs_sel          <= '0';
				Rsrc1_Rscr2_sel   <= '0';
				PC_disable        <= '0';
			END IF;
			IF (opcode = "10100") THEN --JMP
				Flag_Enable       <= '0';
				OutPort_Enable    <= '0';
				RegWrite          <= '0';
				Address           <= '0';
				INT_sig           <= '0';
				MemRead           <= '0';
				MemWrite          <= '0';
				MTR               <= "00";
				SP_sig            <= (others => '0');
				FR                <= '0';
				Write_Data_sel    <= '0';
				RET_sig           <= '0';
				JZ                <= '0';
				JN                <= '0';
				JC                <= '0';
				ALU_sel           <= "000";
				JMP_branch        <= '1';
				UC                <= '1';
				RdRs_sel          <= '0';
				Rsrc1_Rscr2_sel   <= '0';
				PC_disable        <= '0';
			END IF;
			IF (opcode = "10101") THEN --CALL
				Flag_Enable       <= '0';
				OutPort_Enable    <= '0';
				RegWrite          <= '0';
				Address           <= '1';
				INT_sig           <= '0';
				MemRead           <= '0';
				MemWrite          <= '1';
				MTR               <= (others => '0');
				SP_sig            <= "01";
				FR                <= '0';
				Write_Data_sel    <= '1';
				RET_sig           <= '1';
				JZ                <= '0';
				JN                <= '0';
				JC                <= '0';
				ALU_sel           <= "100";
				JMP_branch        <= '1';
				UC                <= '0';
				RdRs_sel          <= '0';
				Rsrc1_Rscr2_sel   <= '0';
				PC_disable        <= '0';
			END IF;
			IF (opcode = "10110") THEN --RET
				Flag_Enable       <= '0';
				OutPort_Enable    <= '0';
				RegWrite          <= '0';
				Address           <= '1';
				INT_sig           <= '0';
				MemRead           <= '1';
				MemWrite          <= '0';
				MTR               <= "01";
				SP_sig            <= "10";
				FR                <= '0';
				Write_Data_sel    <= '0';
				RET_sig           <= '1';
				JZ                <= '0';
				JN                <= '0';
				JC                <= '0';
				ALU_sel           <= "000";
				JMP_branch        <= '1';
				UC                <= '0';
				RdRs_sel          <= '0';
				Rsrc1_Rscr2_sel   <= '0';
				PC_disable        <= '0';
			END IF;
			IF (opcode = "10111") THEN --INT
				Flag_Enable       <= '0';
				OutPort_Enable    <= '0';
				RegWrite          <= '0';
				Address           <= '1';
				INT_sig           <= '1';
				MemRead           <= '0';
				MemWrite          <= '1';
				MTR               <= "00";
				SP_sig            <= "01";
				FR                <= '0';
				Write_Data_sel    <= '1';
				RET_sig           <= '1';
				JZ                <= '0';
				JN                <= '0';
				JC                <= '0';
				ALU_sel           <= "000";
				JMP_branch        <= '1';
				UC                <= '0';
				RdRs_sel          <= '0';
				Rsrc1_Rscr2_sel   <= '0';
				PC_disable        <= '0';
			END IF;
			IF (opcode = "11000") THEN --RTI
				Flag_Enable       <= '0';
				OutPort_Enable    <= '0';
				RegWrite          <= '0';
				Address           <= '1';
				INT_sig           <= '0';
				MemRead           <= '1';
				MemWrite          <= '0';
				MTR               <= "01";
				SP_sig            <= "10";
				FR                <= '1';
				Write_Data_sel    <= '0';
				RET_sig           <= '1';
				JZ                <= '0';
				JN                <= '0';
				JC                <= '0';
				ALU_sel           <= "000";
				JMP_branch        <= '1';
				UC                <= '0';
				RdRs_sel          <= '0';
				Rsrc1_Rscr2_sel   <= '0';
				PC_disable        <= '0';
			END IF;
		END IF;
	END PROCESS;
END Control_Unit_arch;